`include "RegisterFile.sv"
module ID(

);
    
endmodule