`include "../../include/AXI_define.svh"
module Arbiter(
    input clk, rst,
    input 
);
    
endmodule